`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/01/2024 02:02:03 PM
// Design Name: 
// Module Name: InstMem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module InstMem (input [5:0] addr, output [31:0] data_out);
reg [31:0] mem [0:63];
initial begin // Test Program
mem[0] = 32'b00000001010000000000010100010011;
mem[1] = 32'b11111110110000000000010110010011;
mem[2] = 32'b00000010101101010000000001100011;
mem[3] = 32'b00000000101101010001011001100011;
mem[4] = 32'b00000000010100000000101100010011;
mem[5] = 32'b00000000000000000000000001110011;
mem[6] = 32'b00000000101000000000101000010011;
mem[7] = 32'b00000001010001011100100001100011;
mem[8] = 32'b00000000101000000000101110010011;
mem[9] = 32'b00000000000000000000000001110011;
mem[10] = 32'b00000000000100000000111110010011;
mem[11] = 32'b00000000001000000000111100010011;

end
assign data_out = mem[addr];


endmodule